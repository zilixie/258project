module dec_decoder
	(
	input des,
	output [6:0] HEX0, HEX1, HEX2, HEX3
	);
	// Display score in decimal on HEX, every posedge of "des", number
	// increase by 1.
	
	
endmodule