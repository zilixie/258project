module time_control
	(
	input enable,
	output [3:0] plane_amount,
	output [1:0] flying_rate
	);
	// If enable, plane_amount and flying_rate will increase as time pass.
	// plane_amount from 1 to 10, flying_rate from 0 to 3.
	
endmodule